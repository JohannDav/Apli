library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL; 

entity reloj1Hz is  -- ESTE ES EL NOMBRE CORRECTO QUE DEBE USARSE EN TODO EL CÓDIGO
	port (clkin : in STD_LOGIC; -- SEÑAL DE RELOJ DE 50 MHz DEL CRISTAL DE LA TARJETA
											-- CONECTAR AL PIN 12 DE LA EPM240
			clkout : out STD_LOGIC -- SALIDA QUE SERÁ DE 1 Hz (UN PULSO POR SEGUNDO)
);
end reloj1Hz;
architecture funcionamiento of reloj1Hz is
	-- CONTADOR DE 25 BITS: NECESARIO PARA CONTAR HASTA 24,999,999 (25 MILLONES)
	-- 50 MHz / (2 * 1 Hz) - 1 = 24,999,999
	-- CON 25 BITS SE PUEDE CONTAR HASTA 33,554,431 (2^25 - 1)
	signal count: STD_LOGIC_VECTOR ( 24 downto 0 ); -- BIT 24 ES EL MÁS SIGNIFICATIVO (MSB)
													-- BIT 0 ES EL MENOS SIGNIFICATIVO (LSB)
	-- SEÑAL INTERNA TEMPORAL: SE USA PORQUE NO SE PUEDE LEER UNA SALIDA (clkout) 
	-- DENTRO DE UN PROCESS PARA MODIFICARLA
	signal clkint : STD_LOGIC; 
	
	begin
		-- PROCESS: BLOQUE DE CÓDIGO QUE SE EJECUTA SECUENCIALMENTE
		-- SE ACTIVA CADA VEZ QUE LA SEÑAL 'clkin' CAMBIA DE VALOR
		process(clkin)
			begin
				-- DETECTOR DE FLANCO DE SUBIDA: SOLO EJECUTA EL CÓDIGO CUANDO
				-- clkin PASA DE '0' A '1' (DE 0V A 3.3V EN LA TARJETA)
				-- 'event ES UN ATRIBUTO DE VHDL QUE SIGNIFICA "HA OCURRIDO UN EVENTO/CAMBIO"
				if clkin'event and clkin = '1' then 
				
					-- VERIFICA SI EL CONTADOR HA LLEGADO AL VALOR MÁXIMO (24,999,999)
					-- EN BINARIO: "1011111010111100001000000" = 24,999,999 DECIMAL
					if count = "1011111010111100001000000" then 
					
					-- REINICIA EL CONTADOR A CERO (25 BITS EN CERO)
					count <= "0000000000000000000000000";
					
					-- INVIERTE EL VALOR DE clkint: SI ERA '0' PASA A '1', SI ERA '1' PASA A '0'
					-- ESTO OCURRE CADA 25 MILLONES DE CICLOS DE RELOJ = 0.5 SEGUNDOS
					clkint <= not clkint;
					
					-- ASIGNA EL VALOR DE clkint A LA SALIDA clkout
					-- IMPORTANTE: ESTA ASIGNACIÓN ESTÁ DENTRO DEL IF, POR LO QUE SOLO
					-- SE ACTUALIZA CADA 25M CICLOS. SERÍA MEJOR PONERLA FUERA DEL PROCESS
					clkout <= clkint;
					
						else
						-- SI NO HA LLEGADO AL MÁXIMO, INCREMENTA EL CONTADOR EN 1
						-- count + '1': SUMA EL VALOR BINARIO '1' AL VECTOR count
						-- '1' ES UN STD_LOGIC, NO UN INTEGER (POR ESO LAS COMILLAS)
						count <= count + '1';
						
					end if; -- FIN DEL IF INTERNO (verificación del contador)
					
				end if; -- FIN DEL IF EXTERNO (detección de flanco)
				
			end process; -- FIN DEL PROCESS
			
end funcionamiento; -- FIN DE LA ARCHITECTURE