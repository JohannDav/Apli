library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ejercicio_3 is
	Port (A : in std_logic;
			B : in std_logic;
			C : in std_logic;
			D : in std_logic;
			L1 : out std_logic
			L2 : out std_logic);
end ejercicio_3;

architecture arq of ejercicio_3 is
begin
L1 <= A XOR B XOR C XOR D;
L2 <= ((NOT D) AND (NOT C) AND (A XOR B)) OR
      ((NOT B) AND (NOT A) AND (C XOR D)) OR
      (A AND B AND C AND D);